magic
tech sky130A
timestamp 1717310712
<< nwell >>
rect -5 -20 255 225
rect 390 -25 620 225
<< nmos >>
rect 60 -245 95 -185
rect 160 -245 195 -185
rect 485 -245 525 -185
<< pmos >>
rect 60 10 95 70
rect 160 10 195 70
rect 485 10 525 70
<< ndiff >>
rect 15 -195 60 -185
rect 15 -235 20 -195
rect 40 -235 60 -195
rect 15 -245 60 -235
rect 95 -245 160 -185
rect 195 -195 245 -185
rect 195 -235 220 -195
rect 240 -235 245 -195
rect 195 -245 245 -235
rect 435 -245 485 -185
rect 525 -245 580 -185
<< pdiff >>
rect 15 60 60 70
rect 15 20 20 60
rect 40 20 60 60
rect 15 10 60 20
rect 95 10 160 70
rect 195 60 235 70
rect 195 20 210 60
rect 230 20 235 60
rect 195 10 235 20
rect 435 10 485 70
rect 525 10 580 70
<< ndiffc >>
rect 20 -235 40 -195
rect 220 -235 240 -195
<< pdiffc >>
rect 20 20 40 60
rect 210 20 230 60
<< psubdiff >>
rect 60 -320 195 -310
rect 60 -350 85 -320
rect 170 -350 195 -320
rect 60 -360 195 -350
rect 435 -325 580 -310
rect 435 -350 460 -325
rect 555 -350 580 -325
rect 435 -360 580 -350
<< nsubdiff >>
rect 60 185 195 195
rect 60 155 75 185
rect 175 155 195 185
rect 60 145 195 155
rect 450 185 575 200
rect 450 160 465 185
rect 560 160 575 185
rect 450 145 575 160
<< psubdiffcont >>
rect 85 -350 170 -320
rect 460 -350 555 -325
<< nsubdiffcont >>
rect 75 155 175 185
rect 465 160 560 185
<< poly >>
rect 60 70 95 95
rect 160 70 195 95
rect 485 70 525 100
rect 60 -15 95 10
rect 55 -25 95 -15
rect 55 -45 65 -25
rect 85 -45 95 -25
rect 55 -55 95 -45
rect 60 -185 95 -55
rect 160 -85 195 10
rect 150 -95 195 -85
rect 150 -115 160 -95
rect 185 -115 195 -95
rect 150 -125 195 -115
rect 160 -185 195 -125
rect 485 -75 525 10
rect 485 -95 495 -75
rect 515 -95 525 -75
rect 485 -185 525 -95
rect 60 -280 95 -245
rect 160 -280 195 -245
rect 485 -270 525 -245
<< polycont >>
rect 65 -45 85 -25
rect 160 -115 185 -95
rect 495 -95 515 -75
<< locali >>
rect 60 185 195 195
rect 60 155 75 185
rect 175 155 195 185
rect 60 145 195 155
rect 450 190 575 200
rect 450 160 465 190
rect 565 160 575 190
rect 450 145 575 160
rect 110 120 145 145
rect 490 120 510 145
rect 15 90 235 120
rect 15 60 45 90
rect 15 20 20 60
rect 40 20 45 60
rect 15 10 45 20
rect 55 -20 95 -15
rect -205 -25 95 -20
rect -205 -45 65 -25
rect 85 -45 95 -25
rect -205 -50 95 -45
rect 55 -55 95 -50
rect 115 -30 145 70
rect 205 60 235 90
rect 205 20 210 60
rect 230 20 235 60
rect 205 10 235 20
rect 435 100 510 120
rect 435 10 460 100
rect 115 -60 370 -30
rect 340 -70 370 -60
rect 485 -70 525 -65
rect 340 -75 525 -70
rect 150 -90 195 -85
rect -205 -95 195 -90
rect -205 -115 160 -95
rect 185 -115 195 -95
rect 340 -95 495 -75
rect 515 -95 525 -75
rect 340 -100 525 -95
rect 485 -105 525 -100
rect 550 -75 580 70
rect 550 -105 830 -75
rect -205 -120 195 -115
rect 150 -125 195 -120
rect 15 -195 45 -185
rect 15 -235 20 -195
rect 40 -235 45 -195
rect 15 -310 45 -235
rect 215 -195 245 -185
rect 215 -235 220 -195
rect 240 -235 245 -195
rect 215 -245 245 -235
rect 435 -310 470 -185
rect 550 -245 580 -105
rect 15 -320 200 -310
rect 15 -340 85 -320
rect 60 -350 85 -340
rect 170 -340 200 -320
rect 435 -325 580 -310
rect 170 -350 195 -340
rect 60 -360 195 -350
rect 435 -350 460 -325
rect 555 -350 580 -325
rect 435 -360 580 -350
<< viali >>
rect 75 155 175 185
rect 465 185 565 190
rect 465 160 560 185
rect 560 160 565 185
rect 85 -350 170 -320
rect 460 -350 555 -325
<< metal1 >>
rect -195 190 810 200
rect -195 185 465 190
rect -195 155 75 185
rect 175 160 465 185
rect 565 160 810 190
rect 175 155 810 160
rect -195 145 810 155
rect -190 -320 815 -305
rect -190 -350 85 -320
rect 170 -325 815 -320
rect 170 -350 460 -325
rect 555 -350 815 -325
rect -190 -360 815 -350
<< labels >>
rlabel locali -185 -105 -185 -105 1 in2
rlabel metal1 -160 170 -160 170 1 vdd
rlabel metal1 -135 -335 -135 -335 1 vss
rlabel locali -180 -40 -180 -40 1 in1
rlabel locali -180 -105 -180 -105 1 in2
rlabel locali 790 -90 790 -90 1 out
<< end >>
