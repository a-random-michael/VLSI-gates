magic
tech sky130A
timestamp 1717275542
<< nwell >>
rect -5 -20 255 225
<< nmos >>
rect 60 -245 95 -185
rect 160 -245 195 -185
<< pmos >>
rect 60 10 95 70
rect 160 10 195 70
<< ndiff >>
rect 15 -195 60 -185
rect 15 -235 20 -195
rect 40 -235 60 -195
rect 15 -245 60 -235
rect 95 -195 160 -185
rect 95 -235 115 -195
rect 135 -235 160 -195
rect 95 -245 160 -235
rect 195 -195 245 -185
rect 195 -235 220 -195
rect 240 -235 245 -195
rect 195 -245 245 -235
<< pdiff >>
rect 15 60 60 70
rect 15 20 20 60
rect 40 20 60 60
rect 15 10 60 20
rect 95 10 160 70
rect 195 60 235 70
rect 195 20 210 60
rect 230 20 235 60
rect 195 10 235 20
<< ndiffc >>
rect 20 -235 40 -195
rect 115 -235 135 -195
rect 220 -235 240 -195
<< pdiffc >>
rect 20 20 40 60
rect 210 20 230 60
<< psubdiff >>
rect 60 -320 195 -310
rect 60 -350 85 -320
rect 170 -350 195 -320
rect 60 -360 195 -350
<< nsubdiff >>
rect 60 185 195 195
rect 60 155 75 185
rect 175 155 195 185
rect 60 145 195 155
<< psubdiffcont >>
rect 85 -350 170 -320
<< nsubdiffcont >>
rect 75 155 175 185
<< poly >>
rect 60 70 95 95
rect 160 70 195 95
rect 60 -85 95 10
rect 160 -15 195 10
rect 150 -30 195 -15
rect 150 -50 155 -30
rect 180 -50 195 -30
rect 150 -60 195 -50
rect 50 -95 95 -85
rect 50 -115 60 -95
rect 85 -115 95 -95
rect 50 -125 95 -115
rect 60 -185 95 -125
rect 160 -185 195 -60
rect 60 -280 95 -245
rect 160 -280 195 -245
<< polycont >>
rect 155 -50 180 -30
rect 60 -115 85 -95
<< locali >>
rect 60 185 195 195
rect 60 155 75 185
rect 175 155 195 185
rect 60 145 195 155
rect 110 120 145 145
rect 15 90 145 120
rect 15 60 45 90
rect 15 20 20 60
rect 40 20 45 60
rect 15 10 45 20
rect 205 60 235 70
rect 205 20 210 60
rect 230 20 235 60
rect 150 -20 185 -15
rect -60 -30 185 -20
rect -60 -50 155 -30
rect 180 -50 185 -30
rect -60 -55 185 -50
rect 150 -60 185 -55
rect 50 -90 95 -85
rect -60 -95 95 -90
rect -60 -115 60 -95
rect 85 -115 95 -95
rect -60 -120 95 -115
rect 50 -125 95 -120
rect 205 -135 235 20
rect 110 -165 285 -135
rect 15 -195 45 -185
rect 15 -235 20 -195
rect 40 -235 45 -195
rect 15 -310 45 -235
rect 110 -195 145 -165
rect 110 -235 115 -195
rect 135 -235 145 -195
rect 110 -245 145 -235
rect 215 -195 245 -185
rect 215 -235 220 -195
rect 240 -235 245 -195
rect 215 -310 245 -235
rect 15 -320 245 -310
rect 15 -340 85 -320
rect 60 -350 85 -340
rect 170 -340 245 -320
rect 170 -350 195 -340
rect 60 -360 195 -350
<< labels >>
rlabel locali 75 -335 75 -335 1 vss
rlabel locali 70 175 70 175 1 vdd
rlabel locali -50 -105 -50 -105 1 in1
rlabel locali -40 -40 -40 -40 1 in2
rlabel locali 265 -150 265 -150 1 out
<< end >>
