magic
tech sky130A
timestamp 1717311486
<< nwell >>
rect -5 -20 255 225
rect 390 -25 620 225
<< nmos >>
rect 60 -245 95 -185
rect 160 -245 195 -185
rect 485 -245 525 -185
<< pmos >>
rect 60 10 95 70
rect 160 10 195 70
rect 485 10 525 70
<< ndiff >>
rect 15 -195 60 -185
rect 15 -235 20 -195
rect 40 -235 60 -195
rect 15 -245 60 -235
rect 95 -195 160 -185
rect 95 -235 115 -195
rect 135 -235 160 -195
rect 95 -245 160 -235
rect 195 -195 245 -185
rect 195 -235 220 -195
rect 240 -235 245 -195
rect 195 -245 245 -235
rect 435 -195 485 -185
rect 435 -235 440 -195
rect 465 -235 485 -195
rect 435 -245 485 -235
rect 525 -205 580 -185
rect 525 -230 555 -205
rect 575 -230 580 -205
rect 525 -245 580 -230
<< pdiff >>
rect 15 60 60 70
rect 15 20 20 60
rect 40 20 60 60
rect 15 10 60 20
rect 95 10 160 70
rect 195 60 235 70
rect 195 20 210 60
rect 230 20 235 60
rect 195 10 235 20
rect 435 55 485 70
rect 435 20 440 55
rect 460 20 485 55
rect 435 10 485 20
rect 525 55 580 70
rect 525 20 555 55
rect 575 20 580 55
rect 525 10 580 20
<< ndiffc >>
rect 20 -235 40 -195
rect 115 -235 135 -195
rect 220 -235 240 -195
rect 440 -235 465 -195
rect 555 -230 575 -205
<< pdiffc >>
rect 20 20 40 60
rect 210 20 230 60
rect 440 20 460 55
rect 555 20 575 55
<< psubdiff >>
rect 60 -320 195 -310
rect 60 -350 85 -320
rect 170 -350 195 -320
rect 60 -360 195 -350
rect 435 -325 580 -310
rect 435 -350 460 -325
rect 555 -350 580 -325
rect 435 -360 580 -350
<< nsubdiff >>
rect 60 185 195 195
rect 60 155 75 185
rect 175 155 195 185
rect 60 145 195 155
rect 450 185 575 200
rect 450 160 465 185
rect 560 160 575 185
rect 450 145 575 160
<< psubdiffcont >>
rect 85 -350 170 -320
rect 460 -350 555 -325
<< nsubdiffcont >>
rect 75 155 175 185
rect 465 160 560 185
<< poly >>
rect 60 70 95 95
rect 160 70 195 95
rect 485 70 525 100
rect 60 -85 95 10
rect 160 -15 195 10
rect 150 -30 195 -15
rect 150 -50 155 -30
rect 180 -50 195 -30
rect 150 -60 195 -50
rect 50 -95 95 -85
rect 50 -115 60 -95
rect 85 -115 95 -95
rect 50 -125 95 -115
rect 60 -185 95 -125
rect 160 -185 195 -60
rect 485 -75 525 10
rect 485 -95 495 -75
rect 515 -95 525 -75
rect 485 -185 525 -95
rect 60 -280 95 -245
rect 160 -280 195 -245
rect 485 -270 525 -245
<< polycont >>
rect 155 -50 180 -30
rect 60 -115 85 -95
rect 495 -95 515 -75
<< locali >>
rect 60 185 195 195
rect 60 155 75 185
rect 175 155 195 185
rect 60 145 195 155
rect 450 190 575 200
rect 450 160 465 190
rect 565 160 575 190
rect 450 145 575 160
rect 110 120 145 145
rect 490 120 510 145
rect 15 90 145 120
rect 435 100 510 120
rect 15 60 45 90
rect 15 20 20 60
rect 40 20 45 60
rect 15 10 45 20
rect 205 60 235 70
rect 205 20 210 60
rect 230 20 235 60
rect 150 -20 185 -15
rect -200 -30 185 -20
rect -200 -50 155 -30
rect 180 -50 185 -30
rect -200 -55 185 -50
rect 150 -60 185 -55
rect 50 -90 95 -85
rect -205 -95 95 -90
rect -205 -115 60 -95
rect 85 -115 95 -95
rect -205 -120 95 -115
rect 50 -125 95 -120
rect 205 -135 235 20
rect 435 55 465 100
rect 435 20 440 55
rect 460 20 465 55
rect 435 10 465 20
rect 550 55 580 70
rect 550 20 555 55
rect 575 20 580 55
rect 485 -70 525 -65
rect 340 -75 525 -70
rect 340 -95 495 -75
rect 515 -95 525 -75
rect 340 -100 525 -95
rect 340 -135 375 -100
rect 485 -105 525 -100
rect 550 -75 580 20
rect 550 -105 830 -75
rect 110 -165 375 -135
rect 15 -195 45 -185
rect 15 -235 20 -195
rect 40 -235 45 -195
rect 15 -310 45 -235
rect 110 -195 145 -165
rect 110 -235 115 -195
rect 135 -235 145 -195
rect 110 -245 145 -235
rect 215 -195 245 -185
rect 215 -235 220 -195
rect 240 -235 245 -195
rect 215 -310 245 -235
rect 15 -320 245 -310
rect 15 -340 85 -320
rect 60 -350 85 -340
rect 170 -340 245 -320
rect 435 -195 470 -185
rect 435 -235 440 -195
rect 465 -235 470 -195
rect 435 -310 470 -235
rect 550 -205 580 -105
rect 550 -230 555 -205
rect 575 -230 580 -205
rect 550 -245 580 -230
rect 435 -325 580 -310
rect 170 -350 195 -340
rect 60 -360 195 -350
rect 435 -350 460 -325
rect 555 -350 580 -325
rect 435 -360 580 -350
<< viali >>
rect 75 155 175 185
rect 465 185 565 190
rect 465 160 560 185
rect 560 160 565 185
rect 85 -350 170 -320
rect 460 -350 555 -325
<< metal1 >>
rect -195 190 810 200
rect -195 185 465 190
rect -195 155 75 185
rect 175 160 465 185
rect 565 160 810 190
rect 175 155 810 160
rect -195 145 810 155
rect -190 -320 815 -305
rect -190 -350 85 -320
rect 170 -325 815 -320
rect 170 -350 460 -325
rect 555 -350 815 -325
rect -190 -360 815 -350
<< labels >>
rlabel locali -185 -105 -185 -105 1 in2
rlabel metal1 -160 170 -160 170 1 vdd
rlabel metal1 -135 -335 -135 -335 1 vss
rlabel locali 800 -90 800 -90 1 out
rlabel locali -185 -45 -185 -45 1 in1
<< end >>
